module memory_access (
    input clk, rst
);
    
endmodule